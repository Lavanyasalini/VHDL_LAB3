-- write code here
